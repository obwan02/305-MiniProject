library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity game_state_machine is port(Clk: in std_logic);
end entity game_state_machine;

architecture behave of game_state_machine is

begin

end architecture;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pipes is
    port(
        PipeWidth: out signed(9 downto 0);
        PipeHeight: out signed(9 downto 0);
    )
end entity;

architecture construction of pipes is
begin

end architecture;
